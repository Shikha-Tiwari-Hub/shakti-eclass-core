`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif

`ifdef BSV_ASYNC_RESET
 `define BSV_ARESET_EDGE_META or `BSV_RESET_EDGE RST
`else
 `define BSV_ARESET_EDGE_META
`endif

`ifdef BSV_RESET_FIFO_HEAD
 `define BSV_ARESET_EDGE_HEAD `BSV_ARESET_EDGE_META
`else
 `define BSV_ARESET_EDGE_HEAD
`endif

module FIFO2(
   CLK,
   RST,
   D_IN,
   ENQ,
   FULL_N,
   D_OUT,
   DEQ,
   EMPTY_N,
   CLR
);

   parameter width = 1;
   parameter guarded = 1'b1;

   input                     CLK ;
   input                     RST ;
   input [width-1:0]         D_IN;
   input                     ENQ;
   input                     DEQ;
   input                     CLR ;

   output                    FULL_N;
   output                    EMPTY_N;
   output [width-1:0]        D_OUT;

   reg                        full_reg;
   reg                        empty_reg;
   reg [width-1:0]            data0_reg;
   reg [width-1:0]            data1_reg;

   reg                        deqerror;
   reg                        enqerror;

   assign FULL_N = full_reg ;
   assign EMPTY_N = empty_reg ;
   assign D_OUT = data0_reg ;

   wire d0di = (ENQ && !empty_reg) || (ENQ && DEQ && full_reg);
   wire d0d1 = DEQ && !full_reg;
   wire d0h  = ((!DEQ && !ENQ) || (!DEQ && empty_reg) || (!ENQ && full_reg));
   wire d1di = ENQ && empty_reg;

`ifndef BSV_NO_INITIAL_BLOCKS
   // synopsys translate_off
   initial begin
       // Initialize data registers safely
       reg [((width+1)/2)*2-1:0] tmp0, tmp1;
       tmp0 = {((width+1)/2){2'b10}};
       tmp1 = {((width+1)/2){2'b10}};
       data0_reg = tmp0[width-1:0];
       data1_reg = tmp1[width-1:0];

       empty_reg = 1'b0;
       full_reg  = 1'b1;
   end
   // synopsys translate_on
`endif

   // Sequential logic for full/empty registers
   always @(posedge CLK `BSV_ARESET_EDGE_META) begin
      if (RST == `BSV_RESET_VALUE) begin
         empty_reg <= `BSV_ASSIGNMENT_DELAY 1'b0;
         full_reg  <= `BSV_ASSIGNMENT_DELAY 1'b1;
      end else if (CLR) begin
         empty_reg <= `BSV_ASSIGNMENT_DELAY 1'b0;
         full_reg  <= `BSV_ASSIGNMENT_DELAY 1'b1;
      end else if (ENQ && !DEQ) begin
         empty_reg <= `BSV_ASSIGNMENT_DELAY 1'b1;
         full_reg  <= `BSV_ASSIGNMENT_DELAY !empty_reg;
      end else if (DEQ && !ENQ) begin
         full_reg  <= `BSV_ASSIGNMENT_DELAY 1'b1;
         empty_reg <= `BSV_ASSIGNMENT_DELAY !full_reg;
      end
   end

   // Sequential logic for FIFO data registers
   always @(posedge CLK `BSV_ARESET_EDGE_HEAD) begin
`ifdef BSV_RESET_FIFO_HEAD
      if (RST == `BSV_RESET_VALUE) begin
         data0_reg <= `BSV_ASSIGNMENT_DELAY {width{1'b0}};
         data1_reg <= `BSV_ASSIGNMENT_DELAY {width{1'b0}};
      end else
`endif
      begin
         data0_reg <= `BSV_ASSIGNMENT_DELAY
                      ({width{d0di}} & D_IN) |
                      ({width{d0d1}} & data1_reg) |
                      ({width{d0h}} & data0_reg);

         data1_reg <= `BSV_ASSIGNMENT_DELAY
                      d1di ? D_IN : data1_reg;
      end
   end

   // Error checking
   // synopsys translate_off
   always @(posedge CLK) begin
       deqerror = 0;
       enqerror = 0;

       if (RST != `BSV_RESET_VALUE) begin
           if (!empty_reg && DEQ) begin
               deqerror = 1;
               $display("Warning: FIFO2: %m -- Dequeuing from empty fifo");
           end
           if (!full_reg && ENQ && (!DEQ || guarded)) begin
               enqerror = 1;
               $display("Warning: FIFO2: %m -- Enqueuing to a full fifo");
           end
       end
   end
   // synopsys translate_on

endmodule
